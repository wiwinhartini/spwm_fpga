`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 06/21/2022 07:00:39 PM
// Design Name: 
// Module Name: LUT_tap
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module LUT_tbp(
    input clk_in ,
    output reg  [11:0] sine_tbp
    );
parameter SIZE = 407;    // USER INPUT
reg  [11:0] tbp_value [SIZE-1:0];
integer i;

initial begin 
tbp_value[0]=594;
tbp_value[1]=599;
tbp_value[2]=605;
tbp_value[3]=611;
tbp_value[4]=617;
tbp_value[5]=622;
tbp_value[6]=628;
tbp_value[7]=634;
tbp_value[8]=641;
tbp_value[9]=647;
tbp_value[10]=653;
tbp_value[11]=659;
tbp_value[12]=666;
tbp_value[13]=672;
tbp_value[14]=679;
tbp_value[15]=686;
tbp_value[16]=692;
tbp_value[17]=699;
tbp_value[18]=706;
tbp_value[19]=713;
tbp_value[20]=720;
tbp_value[21]=727;
tbp_value[22]=734;
tbp_value[23]=741;
tbp_value[24]=748;
tbp_value[25]=755;
tbp_value[26]=762;
tbp_value[27]=769;
tbp_value[28]=776;
tbp_value[29]=784;
tbp_value[30]=791;
tbp_value[31]=798;
tbp_value[32]=805;
tbp_value[33]=813;
tbp_value[34]=820;
tbp_value[35]=827;
tbp_value[36]=834;
tbp_value[37]=842;
tbp_value[38]=849;
tbp_value[39]=856;
tbp_value[40]=863;
tbp_value[41]=870;
tbp_value[42]=878;
tbp_value[43]=885;
tbp_value[44]=892;
tbp_value[45]=899;
tbp_value[46]=906;
tbp_value[47]=913;
tbp_value[48]=920;
tbp_value[49]=927;
tbp_value[50]=934;
tbp_value[51]=941;
tbp_value[52]=947;
tbp_value[53]=954;
tbp_value[54]=961;
tbp_value[55]=967;
tbp_value[56]=974;
tbp_value[57]=980;
tbp_value[58]=986;
tbp_value[59]=993;
tbp_value[60]=999;
tbp_value[61]=1005;
tbp_value[62]=1011;
tbp_value[63]=1017;
tbp_value[64]=1023;
tbp_value[65]=1029;
tbp_value[66]=1034;
tbp_value[67]=1040;
tbp_value[68]=1045;
tbp_value[69]=1051;
tbp_value[70]=1056;
tbp_value[71]=1061;
tbp_value[72]=1066;
tbp_value[73]=1072;
tbp_value[74]=1076;
tbp_value[75]=1081;
tbp_value[76]=1086;
tbp_value[77]=1091;
tbp_value[78]=1095;
tbp_value[79]=1100;
tbp_value[80]=1104;
tbp_value[81]=1108;
tbp_value[82]=1112;
tbp_value[83]=1116;
tbp_value[84]=1120;
tbp_value[85]=1124;
tbp_value[86]=1128;
tbp_value[87]=1131;
tbp_value[88]=1135;
tbp_value[89]=1138;
tbp_value[90]=1142;
tbp_value[91]=1145;
tbp_value[92]=1148;
tbp_value[93]=1151;
tbp_value[94]=1154;
tbp_value[95]=1157;
tbp_value[96]=1160;
tbp_value[97]=1162;
tbp_value[98]=1165;
tbp_value[99]=1168;
tbp_value[100]=1170;
tbp_value[101]=1172;
tbp_value[102]=1174;
tbp_value[103]=1177;
tbp_value[104]=1179;
tbp_value[105]=1181;
tbp_value[106]=1183;
tbp_value[107]=1184;
tbp_value[108]=1186;
tbp_value[109]=1188;
tbp_value[110]=1189;
tbp_value[111]=1191;
tbp_value[112]=1192;
tbp_value[113]=1194;
tbp_value[114]=1195;
tbp_value[115]=1196;
tbp_value[116]=1198;
tbp_value[117]=1199;
tbp_value[118]=1200;
tbp_value[119]=1201;
tbp_value[120]=1202;
tbp_value[121]=1202;
tbp_value[122]=1203;
tbp_value[123]=1204;
tbp_value[124]=1205;
tbp_value[125]=1205;
tbp_value[126]=1206;
tbp_value[127]=1206;
tbp_value[128]=1207;
tbp_value[129]=1207;
tbp_value[130]=1207;
tbp_value[131]=1208;
tbp_value[132]=1208;
tbp_value[133]=1208;
tbp_value[134]=1208;
tbp_value[135]=1208;
tbp_value[136]=1208;
tbp_value[137]=1208;
tbp_value[138]=1208;
tbp_value[139]=1208;
tbp_value[140]=1208;
tbp_value[141]=1208;
tbp_value[142]=1207;
tbp_value[143]=1207;
tbp_value[144]=1206;
tbp_value[145]=1206;
tbp_value[146]=1205;
tbp_value[147]=1205;
tbp_value[148]=1204;
tbp_value[149]=1203;
tbp_value[150]=1203;
tbp_value[151]=1202;
tbp_value[152]=1201;
tbp_value[153]=1200;
tbp_value[154]=1199;
tbp_value[155]=1198;
tbp_value[156]=1197;
tbp_value[157]=1196;
tbp_value[158]=1194;
tbp_value[159]=1193;
tbp_value[160]=1191;
tbp_value[161]=1190;
tbp_value[162]=1188;
tbp_value[163]=1187;
tbp_value[164]=1185;
tbp_value[165]=1183;
tbp_value[166]=1181;
tbp_value[167]=1179;
tbp_value[168]=1177;
tbp_value[169]=1175;
tbp_value[170]=1173;
tbp_value[171]=1171;
tbp_value[172]=1168;
tbp_value[173]=1166;
tbp_value[174]=1163;
tbp_value[175]=1161;
tbp_value[176]=1158;
tbp_value[177]=1155;
tbp_value[178]=1152;
tbp_value[179]=1149;
tbp_value[180]=1146;
tbp_value[181]=1143;
tbp_value[182]=1140;
tbp_value[183]=1136;
tbp_value[184]=1133;
tbp_value[185]=1129;
tbp_value[186]=1125;
tbp_value[187]=1122;
tbp_value[188]=1118;
tbp_value[189]=1114;
tbp_value[190]=1110;
tbp_value[191]=1105;
tbp_value[192]=1101;
tbp_value[193]=1097;
tbp_value[194]=1092;
tbp_value[195]=1088;
tbp_value[196]=1083;
tbp_value[197]=1078;
tbp_value[198]=1073;
tbp_value[199]=1068;
tbp_value[200]=1063;
tbp_value[201]=1058;
tbp_value[202]=1053;
tbp_value[203]=1047;
tbp_value[204]=1042;
tbp_value[205]=1036;
tbp_value[206]=1031;
tbp_value[207]=1025;
tbp_value[208]=1019;
tbp_value[209]=1013;
tbp_value[210]=1007;
tbp_value[211]=1001;
tbp_value[212]=995;
tbp_value[213]=988;
tbp_value[214]=982;
tbp_value[215]=976;
tbp_value[216]=969;
tbp_value[217]=963;
tbp_value[218]=956;
tbp_value[219]=950;
tbp_value[220]=943;
tbp_value[221]=936;
tbp_value[222]=929;
tbp_value[223]=922;
tbp_value[224]=915;
tbp_value[225]=908;
tbp_value[226]=901;
tbp_value[227]=894;
tbp_value[228]=887;
tbp_value[229]=880;
tbp_value[230]=873;
tbp_value[231]=866;
tbp_value[232]=858;
tbp_value[233]=851;
tbp_value[234]=844;
tbp_value[235]=837;
tbp_value[236]=830;
tbp_value[237]=822;
tbp_value[238]=815;
tbp_value[239]=808;
tbp_value[240]=800;
tbp_value[241]=793;
tbp_value[242]=786;
tbp_value[243]=779;
tbp_value[244]=771;
tbp_value[245]=764;
tbp_value[246]=757;
tbp_value[247]=750;
tbp_value[248]=743;
tbp_value[249]=736;
tbp_value[250]=729;
tbp_value[251]=722;
tbp_value[252]=715;
tbp_value[253]=708;
tbp_value[254]=701;
tbp_value[255]=694;
tbp_value[256]=688;
tbp_value[257]=681;
tbp_value[258]=675;
tbp_value[259]=668;
tbp_value[260]=662;
tbp_value[261]=655;
tbp_value[262]=649;
tbp_value[263]=643;
tbp_value[264]=636;
tbp_value[265]=630;
tbp_value[266]=624;
tbp_value[267]=619;
tbp_value[268]=613;
tbp_value[269]=607;
tbp_value[270]=601;
tbp_value[271]=596;
tbp_value[272]=590;
tbp_value[273]=585;
tbp_value[274]=580;
tbp_value[275]=574;
tbp_value[276]=569;
tbp_value[277]=564;
tbp_value[278]=560;
tbp_value[279]=555;
tbp_value[280]=550;
tbp_value[281]=545;
tbp_value[282]=541;
tbp_value[283]=537;
tbp_value[284]=532;
tbp_value[285]=528;
tbp_value[286]=524;
tbp_value[287]=520;
tbp_value[288]=516;
tbp_value[289]=512;
tbp_value[290]=509;
tbp_value[291]=505;
tbp_value[292]=502;
tbp_value[293]=498;
tbp_value[294]=495;
tbp_value[295]=492;
tbp_value[296]=489;
tbp_value[297]=486;
tbp_value[298]=483;
tbp_value[299]=480;
tbp_value[300]=477;
tbp_value[301]=475;
tbp_value[302]=472;
tbp_value[303]=470;
tbp_value[304]=467;
tbp_value[305]=465;
tbp_value[306]=463;
tbp_value[307]=461;
tbp_value[308]=459;
tbp_value[309]=457;
tbp_value[310]=455;
tbp_value[311]=453;
tbp_value[312]=451;
tbp_value[313]=450;
tbp_value[314]=448;
tbp_value[315]=447;
tbp_value[316]=445;
tbp_value[317]=444;
tbp_value[318]=443;
tbp_value[319]=441;
tbp_value[320]=440;
tbp_value[321]=439;
tbp_value[322]=438;
tbp_value[323]=437;
tbp_value[324]=436;
tbp_value[325]=436;
tbp_value[326]=435;
tbp_value[327]=434;
tbp_value[328]=433;
tbp_value[329]=433;
tbp_value[330]=432;
tbp_value[331]=432;
tbp_value[332]=431;
tbp_value[333]=431;
tbp_value[334]=431;
tbp_value[335]=431;
tbp_value[336]=430;
tbp_value[337]=430;
tbp_value[338]=430;
tbp_value[339]=430;
tbp_value[340]=430;
tbp_value[341]=430;
tbp_value[342]=430;
tbp_value[343]=430;
tbp_value[344]=431;
tbp_value[345]=431;
tbp_value[346]=431;
tbp_value[347]=432;
tbp_value[348]=432;
tbp_value[349]=433;
tbp_value[350]=433;
tbp_value[351]=434;
tbp_value[352]=435;
tbp_value[353]=435;
tbp_value[354]=436;
tbp_value[355]=437;
tbp_value[356]=438;
tbp_value[357]=439;
tbp_value[358]=440;
tbp_value[359]=441;
tbp_value[360]=442;
tbp_value[361]=444;
tbp_value[362]=445;
tbp_value[363]=446;
tbp_value[364]=448;
tbp_value[365]=449;
tbp_value[366]=451;
tbp_value[367]=453;
tbp_value[368]=454;
tbp_value[369]=456;
tbp_value[370]=458;
tbp_value[371]=460;
tbp_value[372]=462;
tbp_value[373]=464;
tbp_value[374]=467;
tbp_value[375]=469;
tbp_value[376]=471;
tbp_value[377]=474;
tbp_value[378]=476;
tbp_value[379]=479;
tbp_value[380]=482;
tbp_value[381]=485;
tbp_value[382]=488;
tbp_value[383]=491;
tbp_value[384]=494;
tbp_value[385]=497;
tbp_value[386]=501;
tbp_value[387]=504;
tbp_value[388]=508;
tbp_value[389]=511;
tbp_value[390]=515;
tbp_value[391]=519;
tbp_value[392]=523;
tbp_value[393]=527;
tbp_value[394]=531;
tbp_value[395]=535;
tbp_value[396]=540;
tbp_value[397]=544;
tbp_value[398]=549;
tbp_value[399]=553;
tbp_value[400]=558;
tbp_value[401]=563;
tbp_value[402]=568;
tbp_value[403]=573;
tbp_value[404]=578;
tbp_value[405]=583;
tbp_value[406]=588;
end 
 
 
 
 

//At every positive edge of the clock, output a sine wave sample.
always@(posedge clk_in)
begin
    sine_tbp = tbp_value[i];
    i = i+ 1;
    if(i == SIZE)
        i = 0;
end
endmodule