`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 06/21/2022 07:00:39 PM
// Design Name: 
// Module Name: LUT_tap
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module LUT_bap(
    input clk_in ,
    output reg [11:0] sine_bap
    );
parameter SIZE = 407;    // USER INPUT
reg [11:0] bap_value [SIZE-1:0];
integer i;

initial begin 
bap_value[0]=410;
bap_value[1]=410;
bap_value[2]=410;
bap_value[3]=410;
bap_value[4]=410;
bap_value[5]=411;
bap_value[6]=411;
bap_value[7]=412;
bap_value[8]=412;
bap_value[9]=413;
bap_value[10]=414;
bap_value[11]=415;
bap_value[12]=416;
bap_value[13]=417;
bap_value[14]=419;
bap_value[15]=420;
bap_value[16]=422;
bap_value[17]=423;
bap_value[18]=425;
bap_value[19]=427;
bap_value[20]=429;
bap_value[21]=431;
bap_value[22]=433;
bap_value[23]=435;
bap_value[24]=437;
bap_value[25]=439;
bap_value[26]=442;
bap_value[27]=444;
bap_value[28]=447;
bap_value[29]=450;
bap_value[30]=453;
bap_value[31]=455;
bap_value[32]=458;
bap_value[33]=462;
bap_value[34]=465;
bap_value[35]=468;
bap_value[36]=471;
bap_value[37]=475;
bap_value[38]=478;
bap_value[39]=482;
bap_value[40]=486;
bap_value[41]=489;
bap_value[42]=493;
bap_value[43]=497;
bap_value[44]=501;
bap_value[45]=505;
bap_value[46]=509;
bap_value[47]=514;
bap_value[48]=518;
bap_value[49]=522;
bap_value[50]=527;
bap_value[51]=531;
bap_value[52]=536;
bap_value[53]=540;
bap_value[54]=545;
bap_value[55]=550;
bap_value[56]=555;
bap_value[57]=560;
bap_value[58]=565;
bap_value[59]=570;
bap_value[60]=575;
bap_value[61]=580;
bap_value[62]=585;
bap_value[63]=590;
bap_value[64]=595;
bap_value[65]=601;
bap_value[66]=606;
bap_value[67]=612;
bap_value[68]=617;
bap_value[69]=623;
bap_value[70]=628;
bap_value[71]=634;
bap_value[72]=639;
bap_value[73]=645;
bap_value[74]=651;
bap_value[75]=657;
bap_value[76]=662;
bap_value[77]=668;
bap_value[78]=674;
bap_value[79]=680;
bap_value[80]=686;
bap_value[81]=692;
bap_value[82]=698;
bap_value[83]=704;
bap_value[84]=710;
bap_value[85]=716;
bap_value[86]=722;
bap_value[87]=728;
bap_value[88]=734;
bap_value[89]=740;
bap_value[90]=746;
bap_value[91]=753;
bap_value[92]=759;
bap_value[93]=765;
bap_value[94]=771;
bap_value[95]=777;
bap_value[96]=783;
bap_value[97]=790;
bap_value[98]=796;
bap_value[99]=802;
bap_value[100]=808;
bap_value[101]=815;
bap_value[102]=821;
bap_value[103]=827;
bap_value[104]=833;
bap_value[105]=839;
bap_value[106]=846;
bap_value[107]=852;
bap_value[108]=858;
bap_value[109]=864;
bap_value[110]=870;
bap_value[111]=877;
bap_value[112]=883;
bap_value[113]=889;
bap_value[114]=895;
bap_value[115]=901;
bap_value[116]=907;
bap_value[117]=913;
bap_value[118]=920;
bap_value[119]=926;
bap_value[120]=932;
bap_value[121]=938;
bap_value[122]=944;
bap_value[123]=950;
bap_value[124]=955;
bap_value[125]=961;
bap_value[126]=967;
bap_value[127]=973;
bap_value[128]=979;
bap_value[129]=985;
bap_value[130]=990;
bap_value[131]=996;
bap_value[132]=1002;
bap_value[133]=1007;
bap_value[134]=1013;
bap_value[135]=1019;
bap_value[136]=1024;
bap_value[137]=1030;
bap_value[138]=1035;
bap_value[139]=1040;
bap_value[140]=1046;
bap_value[141]=1051;
bap_value[142]=1056;
bap_value[143]=1061;
bap_value[144]=1066;
bap_value[145]=1071;
bap_value[146]=1076;
bap_value[147]=1081;
bap_value[148]=1086;
bap_value[149]=1091;
bap_value[150]=1096;
bap_value[151]=1100;
bap_value[152]=1105;
bap_value[153]=1110;
bap_value[154]=1114;
bap_value[155]=1118;
bap_value[156]=1123;
bap_value[157]=1127;
bap_value[158]=1131;
bap_value[159]=1135;
bap_value[160]=1139;
bap_value[161]=1143;
bap_value[162]=1147;
bap_value[163]=1151;
bap_value[164]=1155;
bap_value[165]=1158;
bap_value[166]=1162;
bap_value[167]=1165;
bap_value[168]=1169;
bap_value[169]=1172;
bap_value[170]=1175;
bap_value[171]=1178;
bap_value[172]=1181;
bap_value[173]=1184;
bap_value[174]=1187;
bap_value[175]=1190;
bap_value[176]=1193;
bap_value[177]=1195;
bap_value[178]=1198;
bap_value[179]=1200;
bap_value[180]=1202;
bap_value[181]=1205;
bap_value[182]=1207;
bap_value[183]=1209;
bap_value[184]=1211;
bap_value[185]=1213;
bap_value[186]=1214;
bap_value[187]=1216;
bap_value[188]=1217;
bap_value[189]=1219;
bap_value[190]=1220;
bap_value[191]=1222;
bap_value[192]=1223;
bap_value[193]=1224;
bap_value[194]=1225;
bap_value[195]=1226;
bap_value[196]=1226;
bap_value[197]=1227;
bap_value[198]=1227;
bap_value[199]=1228;
bap_value[200]=1228;
bap_value[201]=1229;
bap_value[202]=1229;
bap_value[203]=1229;
bap_value[204]=1229;
bap_value[205]=1229;
bap_value[206]=1228;
bap_value[207]=1228;
bap_value[208]=1228;
bap_value[209]=1227;
bap_value[210]=1227;
bap_value[211]=1226;
bap_value[212]=1225;
bap_value[213]=1224;
bap_value[214]=1223;
bap_value[215]=1222;
bap_value[216]=1221;
bap_value[217]=1220;
bap_value[218]=1218;
bap_value[219]=1217;
bap_value[220]=1215;
bap_value[221]=1214;
bap_value[222]=1212;
bap_value[223]=1210;
bap_value[224]=1208;
bap_value[225]=1206;
bap_value[226]=1204;
bap_value[227]=1202;
bap_value[228]=1200;
bap_value[229]=1197;
bap_value[230]=1195;
bap_value[231]=1192;
bap_value[232]=1190;
bap_value[233]=1187;
bap_value[234]=1184;
bap_value[235]=1181;
bap_value[236]=1178;
bap_value[237]=1175;
bap_value[238]=1172;
bap_value[239]=1169;
bap_value[240]=1166;
bap_value[241]=1162;
bap_value[242]=1159;
bap_value[243]=1155;
bap_value[244]=1152;
bap_value[245]=1148;
bap_value[246]=1144;
bap_value[247]=1140;
bap_value[248]=1136;
bap_value[249]=1133;
bap_value[250]=1128;
bap_value[251]=1124;
bap_value[252]=1120;
bap_value[253]=1116;
bap_value[254]=1112;
bap_value[255]=1107;
bap_value[256]=1103;
bap_value[257]=1098;
bap_value[258]=1093;
bap_value[259]=1089;
bap_value[260]=1084;
bap_value[261]=1079;
bap_value[262]=1074;
bap_value[263]=1069;
bap_value[264]=1064;
bap_value[265]=1059;
bap_value[266]=1054;
bap_value[267]=1049;
bap_value[268]=1044;
bap_value[269]=1038;
bap_value[270]=1033;
bap_value[271]=1028;
bap_value[272]=1022;
bap_value[273]=1017;
bap_value[274]=1011;
bap_value[275]=1005;
bap_value[276]=1000;
bap_value[277]=994;
bap_value[278]=988;
bap_value[279]=982;
bap_value[280]=977;
bap_value[281]=971;
bap_value[282]=965;
bap_value[283]=959;
bap_value[284]=953;
bap_value[285]=947;
bap_value[286]=941;
bap_value[287]=935;
bap_value[288]=928;
bap_value[289]=922;
bap_value[290]=916;
bap_value[291]=910;
bap_value[292]=904;
bap_value[293]=897;
bap_value[294]=891;
bap_value[295]=885;
bap_value[296]=878;
bap_value[297]=872;
bap_value[298]=866;
bap_value[299]=859;
bap_value[300]=853;
bap_value[301]=846;
bap_value[302]=840;
bap_value[303]=834;
bap_value[304]=827;
bap_value[305]=821;
bap_value[306]=814;
bap_value[307]=808;
bap_value[308]=802;
bap_value[309]=795;
bap_value[310]=789;
bap_value[311]=782;
bap_value[312]=776;
bap_value[313]=770;
bap_value[314]=763;
bap_value[315]=757;
bap_value[316]=751;
bap_value[317]=744;
bap_value[318]=738;
bap_value[319]=732;
bap_value[320]=725;
bap_value[321]=719;
bap_value[322]=713;
bap_value[323]=707;
bap_value[324]=701;
bap_value[325]=695;
bap_value[326]=689;
bap_value[327]=683;
bap_value[328]=677;
bap_value[329]=671;
bap_value[330]=665;
bap_value[331]=659;
bap_value[332]=653;
bap_value[333]=647;
bap_value[334]=642;
bap_value[335]=636;
bap_value[336]=630;
bap_value[337]=625;
bap_value[338]=619;
bap_value[339]=614;
bap_value[340]=608;
bap_value[341]=603;
bap_value[342]=597;
bap_value[343]=592;
bap_value[344]=587;
bap_value[345]=582;
bap_value[346]=577;
bap_value[347]=572;
bap_value[348]=567;
bap_value[349]=562;
bap_value[350]=557;
bap_value[351]=552;
bap_value[352]=547;
bap_value[353]=543;
bap_value[354]=538;
bap_value[355]=534;
bap_value[356]=529;
bap_value[357]=525;
bap_value[358]=520;
bap_value[359]=516;
bap_value[360]=512;
bap_value[361]=508;
bap_value[362]=504;
bap_value[363]=500;
bap_value[364]=496;
bap_value[365]=492;
bap_value[366]=489;
bap_value[367]=485;
bap_value[368]=481;
bap_value[369]=478;
bap_value[370]=474;
bap_value[371]=471;
bap_value[372]=468;
bap_value[373]=465;
bap_value[374]=462;
bap_value[375]=459;
bap_value[376]=456;
bap_value[377]=453;
bap_value[378]=450;
bap_value[379]=448;
bap_value[380]=445;
bap_value[381]=442;
bap_value[382]=440;
bap_value[383]=438;
bap_value[384]=435;
bap_value[385]=433;
bap_value[386]=431;
bap_value[387]=429;
bap_value[388]=427;
bap_value[389]=426;
bap_value[390]=424;
bap_value[391]=422;
bap_value[392]=421;
bap_value[393]=419;
bap_value[394]=418;
bap_value[395]=417;
bap_value[396]=416;
bap_value[397]=415;
bap_value[398]=414;
bap_value[399]=413;
bap_value[400]=412;
bap_value[401]=412;
bap_value[402]=411;
bap_value[403]=411;
bap_value[404]=410;
bap_value[405]=410;
bap_value[406]=410;
end 
 
 

 
//At every positive edge of the clock, output a sine wave sample.
always@(posedge clk_in)
begin
    sine_bap = bap_value[i];
    i = i+ 1;
    if(i == SIZE)
        i = 0;
end
endmodule