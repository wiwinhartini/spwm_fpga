`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 06/21/2022 07:00:39 PM
// Design Name: 
// Module Name: LUT_tap
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module LUT_tap(
    input clk_in ,
    output reg [11:0] sine_tap
    );
parameter SIZE = 407;    // USER INPUT
reg [11:0] tap_value [SIZE-1:0];
integer i;

initial begin 
 tap_value[0]=1208;
tap_value[1]=1208;
tap_value[2]=1208;
tap_value[3]=1208;
tap_value[4]=1208;
tap_value[5]=1208;
tap_value[6]=1207;
tap_value[7]=1207;
tap_value[8]=1207;
tap_value[9]=1206;
tap_value[10]=1206;
tap_value[11]=1205;
tap_value[12]=1204;
tap_value[13]=1204;
tap_value[14]=1203;
tap_value[15]=1202;
tap_value[16]=1201;
tap_value[17]=1200;
tap_value[18]=1199;
tap_value[19]=1198;
tap_value[20]=1197;
tap_value[21]=1196;
tap_value[22]=1195;
tap_value[23]=1193;
tap_value[24]=1192;
tap_value[25]=1190;
tap_value[26]=1189;
tap_value[27]=1187;
tap_value[28]=1186;
tap_value[29]=1184;
tap_value[30]=1182;
tap_value[31]=1180;
tap_value[32]=1178;
tap_value[33]=1176;
tap_value[34]=1174;
tap_value[35]=1171;
tap_value[36]=1169;
tap_value[37]=1167;
tap_value[38]=1164;
tap_value[39]=1162;
tap_value[40]=1159;
tap_value[41]=1156;
tap_value[42]=1153;
tap_value[43]=1150;
tap_value[44]=1147;
tap_value[45]=1144;
tap_value[46]=1141;
tap_value[47]=1137;
tap_value[48]=1134;
tap_value[49]=1130;
tap_value[50]=1127;
tap_value[51]=1123;
tap_value[52]=1119;
tap_value[53]=1115;
tap_value[54]=1111;
tap_value[55]=1107;
tap_value[56]=1103;
tap_value[57]=1098;
tap_value[58]=1094;
tap_value[59]=1089;
tap_value[60]=1084;
tap_value[61]=1080;
tap_value[62]=1075;
tap_value[63]=1070;
tap_value[64]=1065;
tap_value[65]=1060;
tap_value[66]=1054;
tap_value[67]=1049;
tap_value[68]=1044;
tap_value[69]=1038;
tap_value[70]=1032;
tap_value[71]=1027;
tap_value[72]=1021;
tap_value[73]=1015;
tap_value[74]=1009;
tap_value[75]=1003;
tap_value[76]=997;
tap_value[77]=991;
tap_value[78]=984;
tap_value[79]=978;
tap_value[80]=971;
tap_value[81]=965;
tap_value[82]=958;
tap_value[83]=952;
tap_value[84]=945;
tap_value[85]=938;
tap_value[86]=931;
tap_value[87]=925;
tap_value[88]=918;
tap_value[89]=911;
tap_value[90]=904;
tap_value[91]=897;
tap_value[92]=890;
tap_value[93]=882;
tap_value[94]=875;
tap_value[95]=868;
tap_value[96]=861;
tap_value[97]=854;
tap_value[98]=846;
tap_value[99]=839;
tap_value[100]=832;
tap_value[101]=825;
tap_value[102]=817;
tap_value[103]=810;
tap_value[104]=803;
tap_value[105]=796;
tap_value[106]=788;
tap_value[107]=781;
tap_value[108]=774;
tap_value[109]=767;
tap_value[110]=760;
tap_value[111]=752;
tap_value[112]=745;
tap_value[113]=738;
tap_value[114]=731;
tap_value[115]=724;
tap_value[116]=717;
tap_value[117]=710;
tap_value[118]=704;
tap_value[119]=697;
tap_value[120]=690;
tap_value[121]=683;
tap_value[122]=677;
tap_value[123]=670;
tap_value[124]=664;
tap_value[125]=657;
tap_value[126]=651;
tap_value[127]=645;
tap_value[128]=639;
tap_value[129]=632;
tap_value[130]=626;
tap_value[131]=620;
tap_value[132]=615;
tap_value[133]=609;
tap_value[134]=603;
tap_value[135]=598;
tap_value[136]=592;
tap_value[137]=587;
tap_value[138]=581;
tap_value[139]=576;
tap_value[140]=571;
tap_value[141]=566;
tap_value[142]=561;
tap_value[143]=556;
tap_value[144]=552;
tap_value[145]=547;
tap_value[146]=542;
tap_value[147]=538;
tap_value[148]=534;
tap_value[149]=530;
tap_value[150]=525;
tap_value[151]=521;
tap_value[152]=517;
tap_value[153]=514;
tap_value[154]=510;
tap_value[155]=506;
tap_value[156]=503;
tap_value[157]=499;
tap_value[158]=496;
tap_value[159]=493;
tap_value[160]=490;
tap_value[161]=487;
tap_value[162]=484;
tap_value[163]=481;
tap_value[164]=478;
tap_value[165]=476;
tap_value[166]=473;
tap_value[167]=470;
tap_value[168]=468;
tap_value[169]=466;
tap_value[170]=464;
tap_value[171]=461;
tap_value[172]=459;
tap_value[173]=457;
tap_value[174]=456;
tap_value[175]=454;
tap_value[176]=452;
tap_value[177]=450;
tap_value[178]=449;
tap_value[179]=447;
tap_value[180]=446;
tap_value[181]=444;
tap_value[182]=443;
tap_value[183]=442;
tap_value[184]=441;
tap_value[185]=440;
tap_value[186]=439;
tap_value[187]=438;
tap_value[188]=437;
tap_value[189]=436;
tap_value[190]=435;
tap_value[191]=434;
tap_value[192]=434;
tap_value[193]=433;
tap_value[194]=433;
tap_value[195]=432;
tap_value[196]=432;
tap_value[197]=431;
tap_value[198]=431;
tap_value[199]=431;
tap_value[200]=430;
tap_value[201]=430;
tap_value[202]=430;
tap_value[203]=430;
tap_value[204]=430;
tap_value[205]=430;
tap_value[206]=430;
tap_value[207]=430;
tap_value[208]=431;
tap_value[209]=431;
tap_value[210]=431;
tap_value[211]=432;
tap_value[212]=432;
tap_value[213]=433;
tap_value[214]=433;
tap_value[215]=434;
tap_value[216]=434;
tap_value[217]=435;
tap_value[218]=436;
tap_value[219]=437;
tap_value[220]=438;
tap_value[221]=439;
tap_value[222]=440;
tap_value[223]=441;
tap_value[224]=442;
tap_value[225]=443;
tap_value[226]=444;
tap_value[227]=446;
tap_value[228]=447;
tap_value[229]=449;
tap_value[230]=450;
tap_value[231]=452;
tap_value[232]=454;
tap_value[233]=456;
tap_value[234]=457;
tap_value[235]=459;
tap_value[236]=461;
tap_value[237]=464;
tap_value[238]=466;
tap_value[239]=468;
tap_value[240]=470;
tap_value[241]=473;
tap_value[242]=476;
tap_value[243]=478;
tap_value[244]=481;
tap_value[245]=484;
tap_value[246]=487;
tap_value[247]=490;
tap_value[248]=493;
tap_value[249]=496;
tap_value[250]=499;
tap_value[251]=503;
tap_value[252]=506;
tap_value[253]=510;
tap_value[254]=514;
tap_value[255]=517;
tap_value[256]=521;
tap_value[257]=525;
tap_value[258]=530;
tap_value[259]=534;
tap_value[260]=538;
tap_value[261]=542;
tap_value[262]=547;
tap_value[263]=552;
tap_value[264]=556;
tap_value[265]=561;
tap_value[266]=566;
tap_value[267]=571;
tap_value[268]=576;
tap_value[269]=581;
tap_value[270]=587;
tap_value[271]=592;
tap_value[272]=598;
tap_value[273]=603;
tap_value[274]=609;
tap_value[275]=615;
tap_value[276]=620;
tap_value[277]=626;
tap_value[278]=632;
tap_value[279]=639;
tap_value[280]=645;
tap_value[281]=651;
tap_value[282]=657;
tap_value[283]=664;
tap_value[284]=670;
tap_value[285]=677;
tap_value[286]=683;
tap_value[287]=690;
tap_value[288]=697;
tap_value[289]=704;
tap_value[290]=710;
tap_value[291]=717;
tap_value[292]=724;
tap_value[293]=731;
tap_value[294]=738;
tap_value[295]=745;
tap_value[296]=752;
tap_value[297]=760;
tap_value[298]=767;
tap_value[299]=774;
tap_value[300]=781;
tap_value[301]=788;
tap_value[302]=796;
tap_value[303]=803;
tap_value[304]=810;
tap_value[305]=817;
tap_value[306]=825;
tap_value[307]=832;
tap_value[308]=839;
tap_value[309]=846;
tap_value[310]=854;
tap_value[311]=861;
tap_value[312]=868;
tap_value[313]=875;
tap_value[314]=882;
tap_value[315]=890;
tap_value[316]=897;
tap_value[317]=904;
tap_value[318]=911;
tap_value[319]=918;
tap_value[320]=925;
tap_value[321]=931;
tap_value[322]=938;
tap_value[323]=945;
tap_value[324]=952;
tap_value[325]=958;
tap_value[326]=965;
tap_value[327]=971;
tap_value[328]=978;
tap_value[329]=984;
tap_value[330]=991;
tap_value[331]=997;
tap_value[332]=1003;
tap_value[333]=1009;
tap_value[334]=1015;
tap_value[335]=1021;
tap_value[336]=1027;
tap_value[337]=1032;
tap_value[338]=1038;
tap_value[339]=1044;
tap_value[340]=1049;
tap_value[341]=1054;
tap_value[342]=1060;
tap_value[343]=1065;
tap_value[344]=1070;
tap_value[345]=1075;
tap_value[346]=1080;
tap_value[347]=1084;
tap_value[348]=1089;
tap_value[349]=1094;
tap_value[350]=1098;
tap_value[351]=1103;
tap_value[352]=1107;
tap_value[353]=1111;
tap_value[354]=1115;
tap_value[355]=1119;
tap_value[356]=1123;
tap_value[357]=1127;
tap_value[358]=1130;
tap_value[359]=1134;
tap_value[360]=1137;
tap_value[361]=1141;
tap_value[362]=1144;
tap_value[363]=1147;
tap_value[364]=1150;
tap_value[365]=1153;
tap_value[366]=1156;
tap_value[367]=1159;
tap_value[368]=1162;
tap_value[369]=1164;
tap_value[370]=1167;
tap_value[371]=1169;
tap_value[372]=1171;
tap_value[373]=1174;
tap_value[374]=1176;
tap_value[375]=1178;
tap_value[376]=1180;
tap_value[377]=1182;
tap_value[378]=1184;
tap_value[379]=1186;
tap_value[380]=1187;
tap_value[381]=1189;
tap_value[382]=1190;
tap_value[383]=1192;
tap_value[384]=1193;
tap_value[385]=1195;
tap_value[386]=1196;
tap_value[387]=1197;
tap_value[388]=1198;
tap_value[389]=1199;
tap_value[390]=1200;
tap_value[391]=1201;
tap_value[392]=1202;
tap_value[393]=1203;
tap_value[394]=1204;
tap_value[395]=1204;
tap_value[396]=1205;
tap_value[397]=1206;
tap_value[398]=1206;
tap_value[399]=1207;
tap_value[400]=1207;
tap_value[401]=1207;
tap_value[402]=1208;
tap_value[403]=1208;
tap_value[404]=1208;
tap_value[405]=1208;
tap_value[406]=1208;
end 
 


//At every positive edge of the clock, output a sine wave sample.
always@(posedge clk_in)
begin
    sine_tap = tap_value[i];
    i = i+ 1;
    if(i == SIZE)
        i = 0;
end



endmodule